module main
import (
	os
)

fn main () {
	res := os.system("./class_header")
	println(res)
}

