module main

fn main() {
	//hello world
	println('hello')

}
